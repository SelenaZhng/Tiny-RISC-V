//=========================================================================
// 5-Stage Simple Pipelined Processor Datapath
//=========================================================================

`ifndef LAB2_PROC_PROC_ALT_DPATH_V
`define LAB2_PROC_PROC_ALT_DPATH_V

`include "vc/arithmetic.v"
`include "vc/mem-msgs.v"
`include "vc/muxes.v"
`include "vc/regs.v"
`include "vc/regfiles.v"
`include "lab1_imul/IntMulAlt.v"
`include "lab2_proc/tinyrv2_encoding.v"
`include "lab2_proc/ProcDpathImmGen.v"
`include "lab2_proc/ProcDpathAlu.v"

module lab2_proc_ProcAltDpath
#(
  parameter p_num_cores = 1
)
(
  input  logic         clk,
  input  logic         reset,

  // Instruction Memory Port

  output logic [31:0]  imem_reqstream_msg_addr,
  input  mem_resp_4B_t imem_respstream_msg,

  // Data Memory Port

  output logic [31:0]  dmem_reqstream_msg_addr,
  output logic [31:0] dmem_reqstream_msg_data,
  input  logic [31:0]  dmem_respstream_msg_data,

  // mngr communication ports

  input  logic [31:0]  mngr2proc_data,
  output logic [31:0]  proc2mngr_data,

  // control signals (ctrl->dpath)

  input  logic         imem_respstream_drop,

  input  logic         reg_en_F,
  input  logic [1:0]   pc_sel_F,

  input  logic         reg_en_D,
  input  logic         op1_sel_D,
  input  logic [1:0]   op2_sel_D,
  input  logic [1:0]   csrr_sel_D,
  input  logic [2:0]   imm_type_D,
  
  output logic         imul_req_rdy_D,
  input logic          imul_req_val_D,
  input logic  [1:0]   op1_byp_sel_D,
  input logic  [1:0]   op2_byp_sel_D,

  input  logic         reg_en_X,
  input  logic [3:0]   alu_fn_X,
  input  logic [1:0]   ex_result_sel_X,
  
  input logic          imul_resp_rdy_X,
  output logic         imul_resp_val_X,

  input  logic         reg_en_M,
  input  logic         wb_result_sel_M,

  input  logic         reg_en_W,
  input  logic [4:0]   rf_waddr_W,
  input  logic         rf_wen_W,
  input  logic         stats_en_wen_W,

  // status signals (dpath->ctrl)

  output logic [31:0]  inst_D,
  output logic         br_cond_eq_X,
  output logic         br_cond_lt_X,
  output logic         br_cond_ltu_X,

  // extra ports

  input  logic [31:0]  core_id,
  output logic         stats_en
);

  localparam c_reset_vector = 32'h200;
  localparam c_reset_inst   = 32'h00000000;

  // imem addr is just next pc
  assign imem_reqstream_msg_addr = pc_next_F;

  //--------------------------------------------------------------------
  // F stage
  //--------------------------------------------------------------------

  logic [31:0] pc_F;
  logic [31:0] pc_next_F;
  logic [31:0] pc_plus4_F;
  logic [31:0] br_target_X;
  logic [31:0] jal_target_D;
  logic [31:0] jalr_target_X;

  // pc reg (current pc; enable gated by ctrl)
  vc_EnResetReg#(32, c_reset_vector - 32'd4) pc_reg_F
  (
    .clk    (clk),
    .reset  (reset),
    .en     (reg_en_F),
    .d      (pc_next_F),
    .q      (pc_F)
  );

  // pc+4 (sequential next)
  vc_Incrementer#(32, 4) pc_incr_F
  (
    .in   (pc_F),
    .out  (pc_plus4_F)
  );

  logic [31:0] dmem_write_reg_out;
  logic [31:0] alu_result_X;

  // dmem addr/data come from alu + latched rs2
  assign dmem_reqstream_msg_addr = alu_result_X;
  // note: alt path forwards raw alu result (lsb masking handled elsewhere)
  assign jalr_target_X = alu_result_X;
  assign dmem_reqstream_msg_data = dmem_write_reg_out;

  // pc select (seq, branch, jal, jalr)
  vc_Mux4#(32) pc_sel_mux_F
  (
    .in0  (pc_plus4_F),
    .in1  (br_target_X),
    .in2  (jal_target_D),
    .in3  (jalr_target_X),
    .sel  (pc_sel_F),
    .out  (pc_next_F)
  );

  //--------------------------------------------------------------------
  // D stage
  //--------------------------------------------------------------------

  logic [31:0] pc_D;
  logic [ 4:0] inst_rd_D;
  logic [ 4:0] inst_rs1_D;
  logic [ 4:0] inst_rs2_D;
  logic [31:0] imm_D;

  // pipeline pc into D
  vc_EnResetReg#(32) pc_reg_D
  (
    .clk    (clk),
    .reset  (reset),
    .en     (reg_en_D),
    .d      (pc_F),
    .q      (pc_D)
  );

  // pipeline instr into D
  vc_EnResetReg#(32, c_reset_inst) inst_D_reg
  (
    .clk    (clk),
    .reset  (reset),
    .en     (reg_en_D),
    .d      (imem_respstream_msg.data),
    .q      (inst_D)
  );

  // unpack tinyrv2 fields (rs1/rs2/rd etc)
  lab2_proc_tinyrv2_encoding_InstUnpack inst_unpack
  (
    .opcode   (),
    .inst     (inst_D),
    .rs1      (inst_rs1_D),
    .rs2      (inst_rs2_D),
    .rd       (inst_rd_D),
    .funct3   (),
    .funct7   (),
    .csr      ()
  );

  // immediate generator (i/s/b/u/j)
  lab2_proc_ProcDpathImmGen imm_gen_D
  (
    .imm_type (imm_type_D),
    .inst     (inst_D),
    .imm      (imm_D)
  );

  logic [31:0] rf_rdata0_D;
  logic [31:0] rf_rdata1_D;
  logic [31:0] rf_wdata_W;

  // regfile 2r1w, x0 hardwired to zero
  vc_Regfile_2r1w_zero rf
  (
    .clk      (clk),
    .reset    (reset),
    .rd_addr0 (inst_rs1_D),
    .rd_data0 (rf_rdata0_D),
    .rd_addr1 (inst_rs2_D),
    .rd_data1 (rf_rdata1_D),
    .wr_en    (rf_wen_W),
    .wr_addr  (rf_waddr_W),
    .wr_data  (rf_wdata_W)
  );

  logic [31:0] csrr_data_D;
  logic [31:0] num_cores;
  assign num_cores = p_num_cores;

  // csr source select (manager/numcores/coreid)
  vc_Mux3#(32) csrr_sel_mux_D
  (
   .in0  (mngr2proc_data),
   .in1  (num_cores),
   .in2  (core_id),
   .sel  (csrr_sel_D),
   .out  (csrr_data_D)
  );

  logic [31:0] op2_D;

  // op2 select (byp/imm/csr)
  vc_Mux3#(32) op2_sel_mux_D
  (
    .in0  (op2_byp_out_D),
    .in1  (imm_D),
    .in2  (csrr_data_D),
    .sel  (op2_sel_D),
    .out  (op2_D)
  );

  // jal target = pc + imm
  vc_Adder#(32) pc_plus_imm_D
  (
    .in0  (pc_D),
    .in1  (imm_D),
    .cin  (1'b0),
    .out  (jal_target_D),
    .cout ()
  );

  logic [31:0] pc_reg_X_out;

  // pipeline pc into X (for pc+4 calc)
  vc_EnResetReg#(32) pc_reg_X
  (
    .clk   (clk),
    .reset (reset),
    .en    (reg_en_X),
    .d     (pc_D),
    .q     (pc_reg_X_out)
  );

  logic [31:0] op1_sel_mux_out;

  // op1 select (pc vs bypassed rs1)
  vc_Mux2#(32) op1_sel_mux_D
  (
    .in0  (pc_D),
    .in1  (op1_byp_out_D),
    .sel  (op1_sel_D),
    .out  (op1_sel_mux_out)
  );

  // BYPASS MUXES

  logic [31:0] bypass_from_X;
  logic [31:0] bypass_from_M;
  logic [31:0] bypass_from_W;
  logic [31:0] op1_byp_out_D;
  logic [31:0] op2_byp_out_D;

  // op1 bypass pick (W/M/X/rf)
  vc_Mux4#(32) op1_byp_mux_D
  (
    .in0  (bypass_from_W),
    .in1  (bypass_from_M),
    .in2  (bypass_from_X),
    .in3  (rf_rdata0_D),
    .sel  (op1_byp_sel_D),
    .out  (op1_byp_out_D)
  );

  // op2 bypass pick (rf/W/M/X)
  vc_Mux4#(32) op2_byp_mux_D
  (
    .in0  (rf_rdata1_D),
    .in1  (bypass_from_W),
    .in2  (bypass_from_M),
    .in3  (bypass_from_X),
    .sel  (op2_byp_sel_D),
    .out  (op2_byp_out_D)
  );

  //--------------------------------------------------------------------
  // X stage
  //--------------------------------------------------------------------

  logic [31:0] op1_X;
  logic [31:0] op2_X;

  // pipeline alu operands into X
  vc_EnResetReg#(32, 0) op1_reg_X
  (
    .clk   (clk),
    .reset (reset),
    .en    (reg_en_X),
    .d     (op1_sel_mux_out),
    .q     (op1_X)
  );

  vc_EnResetReg#(32, 0) op2_reg_X
  (
    .clk   (clk),
    .reset (reset),
    .en    (reg_en_X),
    .d     (op2_D),
    .q     (op2_X)
  );

  // branch target pipeline reg (pc+imm carried into X)
  vc_EnResetReg#(32, 0) br_target_reg_X
  (
    .clk   (clk),
    .reset (reset),
    .en    (reg_en_X),
    .d     (jal_target_D),
    .q     (br_target_X)
  );

  logic [31:0] ex_result_X;

  // main alu (also spits out compare flags)
  lab2_proc_ProcDpathAlu alu
  (
    .in0      (op1_X),
    .in1      (op2_X),
    .fn       (alu_fn_X),
    .out      (alu_result_X),
    .ops_eq   (br_cond_eq_X),
    .ops_lt   (br_cond_lt_X),
    .ops_ltu  (br_cond_ltu_X)
  );

  logic [31:0] pc_X;
  logic [31:0] imul_resp_msg;

  // select exe result: pc+4 vs alu vs imul
  assign bypass_from_X = ex_result_X;
  vc_Mux3#(32) ex_result_sel_mux_X
  (
    .in0    (pc_X),
    .in1    (alu_result_X),
    .in2    (imul_resp_msg),
    .sel    (ex_result_sel_X),
    .out    (ex_result_X)
  );

  // store data latch (rs2 after bypassing)
  vc_EnResetReg#(32, 0) dmem_write_data_reg_X
  (
    .clk   (clk),
    .reset (reset),
    .en    (reg_en_X),
    .d     (op2_byp_out_D),
    .q     (dmem_write_reg_out)
  );

  // pc+4 in X (for jal writeback)
  vc_Incrementer#(32, 4) pc_incr_X
  (
    .in   (pc_reg_X_out),
    .out  (pc_X)
  );
  
  logic [63:0] imul_req_msg;
  assign imul_req_msg = {op1_sel_mux_out, op2_D};
  
  // iterative int multiplier (req/resp handshake)
  lab1_imul_IntMulAlt imul
  (
    .clk(clk),
    .reset(reset),
    .istream_val(imul_req_val_D),
    .istream_rdy(imul_req_rdy_D),
    .istream_msg(imul_req_msg),
    .ostream_val(imul_resp_val_X),
    .ostream_rdy(imul_resp_rdy_X),
    .ostream_msg(imul_resp_msg) 
  );

  //--------------------------------------------------------------------
  // M stage
  //--------------------------------------------------------------------

  logic [31:0] ex_result_M;

  // pipeline exe result to M
  vc_EnResetReg#(32, 0) ex_result_reg_M
  (
    .clk    (clk),
    .reset  (reset),
    .en     (reg_en_M),
    .d      (ex_result_X),
    .q      (ex_result_M)
  );

  logic [31:0] dmem_result_M;
  logic [31:0] wb_result_M;

  // load data from dmem response
  assign dmem_result_M = dmem_respstream_msg_data;
  // expose M result to bypass net
  assign bypass_from_M = wb_result_M;

  // choose wb source in M (alu/pc vs load)
  vc_Mux2#(32) wb_result_sel_mux_M
  (
    .in0    (ex_result_M),
    .in1    (dmem_result_M),
    .sel    (wb_result_sel_M),
    .out    (wb_result_M)
  );

  //--------------------------------------------------------------------
  // W stage
  //--------------------------------------------------------------------

  logic [31:0] wb_result_W;

  // expose W result to bypass net
  assign bypass_from_W = wb_result_W;

  // pipeline to W (final wb data)
  vc_EnResetReg#(32, 0) wb_result_reg_W
  (
    .clk    (clk),
    .reset  (reset),
    .en     (reg_en_W),
    .d      (wb_result_M),
    .q      (wb_result_W)
  );

  logic [31:0] stats_en_W;
  assign stats_en = | stats_en_W;
  assign proc2mngr_data = wb_result_W;
  assign rf_wdata_W = wb_result_W;

  // stats enable (counts when non-zero in W)
  vc_EnResetReg#(32, 0) stats_en_reg_W
  (
   .clk    (clk),
   .reset  (reset),
   .en     (stats_en_wen_W),
   .d      (wb_result_W),
   .q      (stats_en_W)
  );

endmodule

`endif /* LAB2_PROC_PROC_ALT_DPATH_V */
